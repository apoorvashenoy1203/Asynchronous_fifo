 `define DATA_SIZE 8
`define ADDR_SIZE 4

 package pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "defines.sv"
  `include "fifo_seq_item.sv"
  `include "sequencer.sv"
  `include "sequence.sv"
  `include "write_driver.sv"
  `include "write_monitor.sv"
  `include "read_driver.sv"
  `include "read_monitor.sv"
  `include "fifo_agent.sv"
  `include "fifo_scoreboard.sv"
  `include "subscriber.sv"
  `include "fifo_env.sv"
  `include "test.sv"
endpackage
